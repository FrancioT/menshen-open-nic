
`timescale 1ns / 1ps

module tb_rmt_wrapper_stages #(
    // Slave AXI parameters
	parameter C_S_AXI_DATA_WIDTH = 32,
	parameter C_S_AXI_ADDR_WIDTH = 12,
	parameter C_BASEADDR = 32'h80000000,
	// AXI Stream parameters
	// Slave
	parameter C_S_AXIS_DATA_WIDTH = 512,
	parameter C_S_AXIS_TUSER_WIDTH = 128,
	// Master
	parameter C_M_AXIS_DATA_WIDTH = 512,
	// self-defined
	parameter PHV_ADDR_WIDTH = 4
)();

reg                                 clk;
reg                                 aresetn;

reg [C_S_AXIS_DATA_WIDTH-1:0]		s_axis_tdata;
reg [((C_S_AXIS_DATA_WIDTH/8))-1:0]	s_axis_tkeep;
reg [C_S_AXIS_TUSER_WIDTH-1:0]		s_axis_tuser;
reg									s_axis_tvalid;
wire								s_axis_tready;
reg									s_axis_tlast;

wire [C_S_AXIS_DATA_WIDTH-1:0]		    m_axis_tdata;
wire [((C_S_AXIS_DATA_WIDTH/8))-1:0]    m_axis_tkeep;
wire [C_S_AXIS_TUSER_WIDTH-1:0]		    m_axis_tuser;
wire								    m_axis_tvalid;
reg										m_axis_tready;
wire									m_axis_tlast;


//clk signal
localparam CYCLE = 10;

always begin
    #(CYCLE/2) clk = ~clk;
end

//reset signal
initial begin
    clk = 0;
    aresetn = 1;
    #(10);
    aresetn = 0; //reset all the values
    #(10);
    aresetn = 1;
end


initial begin
	#(3*CYCLE+CYCLE/2);
    #(40* CYCLE)
    m_axis_tready <= 1'b1;
    s_axis_tdata <= 512'b0; 
    s_axis_tkeep <= 64'h0;
    s_axis_tuser <= 128'h0;
    s_axis_tvalid <= 1'b0;
    s_axis_tlast <= 1'b0;

	#(30*CYCLE)
	// conf1.txt:
	s_axis_tdata <= 512'h000000000000000000000000000000010000902f2e00f2f1d204dededede6f6f6f6f0ede1140000001004200004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000270e250d230c910ba108;
	s_axis_tkeep <= 64'h00000000000fffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010005902a2e00f2f1d204dededede6f6f6f6f0ede1140000001004200004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000270e250d230c910ba108;
	s_axis_tkeep <= 64'h00000000000fffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000100014f5e1f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c0000;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f0117ea3300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffff0000ffffffffffffffffffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000275683400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000a00100000000000000000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000f02282d6900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007409c0200001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000001000245683400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000d00000000000000000000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f02292c6900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007409c0100001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010009cf541f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c8001;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f0917e23300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000a35603400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e00100000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000f0ae8246900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007809c0200001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000001000af55d3400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200300000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f0ae9236900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007809c0100001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010011cf4c1f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c8001;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f1117da3300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000001285583400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000900100000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000f12281d6900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007409c0200001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010012a5553400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000700300000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f12291c6900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007409c0100001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010019cf441f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c8001;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f1917d23300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000001a25513400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000f1ae8146900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007809c0200001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000001001a054d3400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100400000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f1ae9136900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007809c0100001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010021cf3c1f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c8001;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f2117ca3300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000002275493400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a00000000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000f22280d6900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007409c0200001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010022b5443400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000600400000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f22290c6900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c003008007409c0100001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)


	// confsys.txt:
	s_axis_tdata <= 512'h0000000000000000000000000000000100214f3e1f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c0000;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f2117ca3300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000200214f3d1f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c0000;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000020f2117c93300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000300214f3c1f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c0000;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000030f2117c83300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000400214f3b1f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c0000;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000040f2117c73300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000f00214f301f00f2f1d204dededede6f6f6f6f1dde1140000001003300004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c0000;
	s_axis_tkeep <= 64'h000000000000001f;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000f0f2117bc3300f2f1d204dededede6f6f6f6f09de1140000001004700004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000080ffffffffffffffff00000000ffffffffffffffffffffffff;
	s_axis_tkeep <= 64'h0000000001ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000002275493400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a00000000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000000f2286596900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000050c50000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000001002265483400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a00000000000000000000000000000002000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000010f2286586900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000050c50000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000002002255473400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a00000000000000000000000000000003000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000020f2286576900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000050c50000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000003002245463400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a00000000000000000000000000000004000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000030f2286566900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000050c50000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000004002295443400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a0000000000000000000000000000000f000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000040f2286556900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000050c50000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000005002285443400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000900000000000000000000000000000001000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000050f228b646900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040c00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000006002275433400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000900000000000000000000000000000002000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000060f228b636900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040c00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000007002265423400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000900000000000000000000000000000003000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000070f228b626900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040c00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000008002255413400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000900000000000000000000000000000004000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000080f228b616900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040c00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000090022a53f3400f2f1d204dededede6f6f6f6f08de1140000001004800004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000090000000000000000000000000000000f000;
	s_axis_tkeep <= 64'h0000000003ffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h000000000000000000000000000000090f228b606900f2f1d204dededede6f6f6f6fd3dd1140000001007d00004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f00000e00100c00300800700000f00001e00003c0000780000f0;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040c00000e00100c00300800700;
	s_axis_tkeep <= 64'h0000000000007fff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)


	// stateconf.txt:
	s_axis_tdata <= 512'h00000000000000000000000000000001001355541c00f2f1d204dededede6f6f6f6f20de1140000001003000004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004;
	s_axis_tkeep <= 64'h0000000000000003;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000002001351531c00f2f1d204dededede6f6f6f6f20de1140000001003000004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000404;
	s_axis_tkeep <= 64'h0000000000000003;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h0000000000000000000000000000000300134d521c00f2f1d204dededede6f6f6f6f20de1140000001003000004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000804;
	s_axis_tkeep <= 64'h0000000000000003;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000004001349511c00f2f1d204dededede6f6f6f6f20de1140000001003000004500080f0000810504030201000b0a09080706;
	s_axis_tkeep <= 64'hffffffffffffffff;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b0;
	#(CYCLE)
	s_axis_tdata <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c04;
	s_axis_tkeep <= 64'h0000000000000003;
	s_axis_tvalid <= 1'b1;
	s_axis_tlast <= 1'b1;
	#CYCLE
	s_axis_tvalid <= 1'b0;
	s_axis_tlast <= 1'b0;
	#(30*CYCLE)


    // test packet
    // padding: 00000000 bit
    // res    : 82000000 = 40 	
    // op_a   : a0000000 = 10
    // op_b   : 50000000 = 5
    // op     : 1a00 = - / 0d00 = +
    //s_axis_tdata <= 512'h0000000026000000050000000a0000000d004c4d1a00e110d204dededede6f6f6f6f22de1140000001002e000045000801000081050403020100090000000000;	
    s_axis_tdata <= 512'h0000000028000000050000000a0000000d004c4d1a00e110d204dededede6f6f6f6f22de1140000001002e000045000801000081050403020100090000000000;	
    s_axis_tkeep <= 64'hffffffffffffffff;
    s_axis_tvalid <= 1'b1;
    s_axis_tlast <= 1'b1;
    #CYCLE
    s_axis_tvalid <= 1'b0;
    s_axis_tlast <= 1'b0;
    
    // Check result
	@(m_axis_tvalid == 1'b1)
	assert (m_axis_tdata[479:472] == 8'h46) $display ("TEST PASSED");
	$finish;
end


rmt_wrapper #(
	.C_S_AXI_DATA_WIDTH(),
	.C_S_AXI_ADDR_WIDTH(),
	.C_BASEADDR(),
	.C_S_AXIS_DATA_WIDTH(C_S_AXIS_DATA_WIDTH),
	.C_S_AXIS_TUSER_WIDTH(),
	.C_M_AXIS_DATA_WIDTH(C_M_AXIS_DATA_WIDTH),
	.PHV_ADDR_WIDTH()
)rmt_wrapper_ins
(
	.clk(clk),		// axis clk
	.aresetn(aresetn),	

	// input Slave AXI Stream
	.s_axis_tdata(s_axis_tdata),
	.s_axis_tkeep(s_axis_tkeep),
	.s_axis_tuser(s_axis_tuser),
	.s_axis_tvalid(s_axis_tvalid),
	.s_axis_tready(s_axis_tready),
	.s_axis_tlast(s_axis_tlast),

	// output Master AXI Stream
	.m_axis_tdata(m_axis_tdata),
	.m_axis_tkeep(m_axis_tkeep),
	.m_axis_tuser(m_axis_tuser),
	.m_axis_tvalid(m_axis_tvalid),
	.m_axis_tready(m_axis_tready),
	.m_axis_tlast(m_axis_tlast)
	
);

endmodule
